module tfgrid

struct Ipaddr {
	// check what we have in crystallib, can prob re-use
}

struct Ipaddr6 {
	// check what we have in crystallib, can prob re-use
}

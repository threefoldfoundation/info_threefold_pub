module tfgrid

// see https://github.com/threefoldtech/zos/tree/zos3/new-types/pkg/gridtypes/zos
